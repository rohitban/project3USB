//Your testbench module
module test
  (output logic clk, rst_L);

  //Set up clk, rst_L, and then call your usbHost.sv tasks here  

  //Ex: host.prelabRequest(data);
  //    host.writeData(memPage, data, success);
  //    host.readData(memPage, data, success);  
    

endmodule
