module bs_encoder

endmodule: bs_encoder
